module mux2x1_1bit(output result, input a, input b, input sel);

	
	


endmodule