module mod_cu(output wire mod_result, input wire clk, input wire start, input[31:0] A, input[31:0} B);

reg curr_state, next_state;

endmodule